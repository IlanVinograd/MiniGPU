`timescale 1ns/1ps

module resp_packet_tx #(

)(
    
);

    
endmodule