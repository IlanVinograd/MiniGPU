`timescale 1ns/1ps

module cmd_status #(
  
)(

);
  
endmodule